--libraries to be used are specified here
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

--entity declaration with port definitions
entity syn_count4 is
port ( clk:     in std_logic;
	reset: in std_logic;
          counter : out std_logic_vector(3 downto 0)
);
end syn_count4;

--architecture of entity
architecture Behavioral of syn_count4 is
--signal declaration.
signal J3,J4,Q1,Q2,Q3,Q4,Qbar1,Qbar2,Qbar3,Qbar4: std_logic :='0';

begin 
J3 <= Q1 and Q2;
J4<= J3 and Q3;

--entity instantiations
FF1 : entity work.JK_Flipflop port map (clk,'1','1',Q1,Qbar1,reset);
FF2 : entity work.JK_Flipflop port map (clk,Q1,Q1,Q2,Qbar2,reset);
FF3 : entity work.JK_Flipflop port map (clk,J3,J3,Q3,Qbar3,reset);
FF4 : entity work.JK_Flipflop port map (clk,J4,J4,Q4,Qbar4,reset);
counter <= Q4 & Q3 & Q2 & Q1;

end Behavioral;